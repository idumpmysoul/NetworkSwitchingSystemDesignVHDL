library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity switch is --only 1 port receiver, 3 port sending
    port (
        fa01    :   inout std_logic_vector(7 downto 0);
        fa02    :   inout 
        fa03

    );
end entity switch;

architecture rtl of switch is
    
begin
    
    
    
end architecture rtl;