library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity EndROM is
    port (
        3
        
    );
end entity EndROM;

architecture rtl of EndROM is
    component register8bit is
        port (
            
        );
    end component register8bit;
begin
    
    
    
end architecture rtl;
