library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity switchport is
    port (
        fa01        : inout std_logic_vector(127 downto 0);
        fa01_add    : inout std_logic_vector(47 downto 0);
        fa02        : inout std_logic_vector(127 downto 0);
        fa02_add    : inout std_logic_vector(47 downto 0);
        fa03        : inout std_logic_vector(127 downto 0);
        fa03_add    : inout std_logic_vector(47 downto 0);
        fa04        : inout std_logic_vector(127 downto 0);
        fa04_add    : inout std_logic_vector(47 downto 0);
        fa05        : inout std_logic_vector(127 downto 0);
        fa05_add    : inout std_logic_vector(47 downto 0);
        fa06        : inout std_logic_vector(127 downto 0);
        fa06_add    : inout std_logic_vector(47 downto 0);
        fa07        : inout std_logic_vector(127 downto 0);
        fa07_add    : inout std_logic_vector(47 downto 0);
        fa08        : inout std_logic_vector(127 downto 0);
        fa08_add    : inout std_logic_vector(47 downto 0);
        fa09        : inout std_logic_vector(127 downto 0);
        fa09_add    : inout std_logic_vector(47 downto 0);
        fa010        : inout std_logic_vector(127 downto 0);
        fa010_add    : inout std_logic_vector(47 downto 0);
        fa011        : inout std_logic_vector(127 downto 0);
        fa011_add    : inout std_logic_vector(47 downto 0);
        fa012        : inout std_logic_vector(127 downto 0);
        fa012_add    : inout std_logic_vector(47 downto 0);
    );
end entity switchport;

architecture rtl of switchport is
    
begin
    
    
    
end architecture rtl;