library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity register8bit is
    port (
        
    );
end entity register8bit;

architecture rtl of register8bit is
    
begin
    
    
    
end architecture rtl;

