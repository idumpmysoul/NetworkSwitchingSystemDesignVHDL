library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity endDevice is
    port (
        mac_add                                                                                                                                                                                                                                                                                                                                                                                                                                  a 
    );
end entity endDevice;

architecture rtl of endDevice is
    
begin
    
    
    
end architecture rtl;