library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity endDevice is
    port (
        frame_in     : 
    );
end entity endDevice;

architecture rtl of endDevice is
    
begin
    
    
    
end architecture rtl;