library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity switch is
    port (
        INPUT   :   in std_logic_vector(7 downto 0);

    );
end entity switch;

architecture rtl of switch is
    
begin
    
    
    
end architecture rtl;